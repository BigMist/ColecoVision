library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d8dfc287",
    12 => x"86c0c84e",
    13 => x"49d8dfc2",
    14 => x"48cccdc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087dfdc",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d60299",
    50 => x"c348d4ff",
    51 => x"526878ff",
    52 => x"484966c4",
    53 => x"a6c888c1",
    54 => x"05997158",
    55 => x"4f2687ea",
    56 => x"ff1e731e",
    57 => x"ffc34bd4",
    58 => x"c34a6b7b",
    59 => x"496b7bff",
    60 => x"b17232c8",
    61 => x"6b7bffc3",
    62 => x"7131c84a",
    63 => x"7bffc3b2",
    64 => x"32c8496b",
    65 => x"4871b172",
    66 => x"4d2687c4",
    67 => x"4b264c26",
    68 => x"5e0e4f26",
    69 => x"0e5d5c5b",
    70 => x"d4ff4a71",
    71 => x"c348724c",
    72 => x"7c7098ff",
    73 => x"bfcccdc2",
    74 => x"d087c805",
    75 => x"30c94866",
    76 => x"d058a6d4",
    77 => x"29d84966",
    78 => x"ffc34871",
    79 => x"d07c7098",
    80 => x"29d04966",
    81 => x"ffc34871",
    82 => x"d07c7098",
    83 => x"29c84966",
    84 => x"ffc34871",
    85 => x"d07c7098",
    86 => x"ffc34866",
    87 => x"727c7098",
    88 => x"7129d049",
    89 => x"98ffc348",
    90 => x"4b6c7c70",
    91 => x"4dfff0c9",
    92 => x"05abffc3",
    93 => x"ffc387d0",
    94 => x"c14b6c7c",
    95 => x"87c6028d",
    96 => x"02abffc3",
    97 => x"487387f0",
    98 => x"1e87fffd",
    99 => x"d4ff49c0",
   100 => x"78ffc348",
   101 => x"c8c381c1",
   102 => x"f104a9b7",
   103 => x"1e4f2687",
   104 => x"87e71e73",
   105 => x"4bdff8c4",
   106 => x"ffc01ec0",
   107 => x"49f7c1f0",
   108 => x"c487dffd",
   109 => x"05a8c186",
   110 => x"ff87eac0",
   111 => x"ffc348d4",
   112 => x"c0c0c178",
   113 => x"1ec0c0c0",
   114 => x"c1f0e1c0",
   115 => x"c1fd49e9",
   116 => x"7086c487",
   117 => x"87ca0598",
   118 => x"c348d4ff",
   119 => x"48c178ff",
   120 => x"e6fe87cb",
   121 => x"058bc187",
   122 => x"c087fdfe",
   123 => x"87defc48",
   124 => x"ff1e731e",
   125 => x"ffc348d4",
   126 => x"c04bd378",
   127 => x"f0ffc01e",
   128 => x"fc49c1c1",
   129 => x"86c487cc",
   130 => x"ca059870",
   131 => x"48d4ff87",
   132 => x"c178ffc3",
   133 => x"fd87cb48",
   134 => x"8bc187f1",
   135 => x"87dbff05",
   136 => x"e9fb48c0",
   137 => x"5b5e0e87",
   138 => x"d4ff0e5c",
   139 => x"87dbfd4c",
   140 => x"c01eeac6",
   141 => x"c8c1f0e1",
   142 => x"87d6fb49",
   143 => x"a8c186c4",
   144 => x"fe87c802",
   145 => x"48c087ea",
   146 => x"fa87e2c1",
   147 => x"497087d2",
   148 => x"99ffffcf",
   149 => x"02a9eac6",
   150 => x"d3fe87c8",
   151 => x"c148c087",
   152 => x"ffc387cb",
   153 => x"4bf1c07c",
   154 => x"7087f4fc",
   155 => x"ebc00298",
   156 => x"c01ec087",
   157 => x"fac1f0ff",
   158 => x"87d6fa49",
   159 => x"987086c4",
   160 => x"c387d905",
   161 => x"496c7cff",
   162 => x"7c7cffc3",
   163 => x"c0c17c7c",
   164 => x"87c40299",
   165 => x"87d548c1",
   166 => x"87d148c0",
   167 => x"c405abc2",
   168 => x"c848c087",
   169 => x"058bc187",
   170 => x"c087fdfe",
   171 => x"87dcf948",
   172 => x"c21e731e",
   173 => x"c148cccd",
   174 => x"ff4bc778",
   175 => x"78c248d0",
   176 => x"ff87c8fb",
   177 => x"78c348d0",
   178 => x"e5c01ec0",
   179 => x"49c0c1d0",
   180 => x"c487fff8",
   181 => x"05a8c186",
   182 => x"c24b87c1",
   183 => x"87c505ab",
   184 => x"f9c048c0",
   185 => x"058bc187",
   186 => x"fc87d0ff",
   187 => x"cdc287f7",
   188 => x"987058d0",
   189 => x"c187cd05",
   190 => x"f0ffc01e",
   191 => x"f849d0c1",
   192 => x"86c487d0",
   193 => x"c348d4ff",
   194 => x"fdc278ff",
   195 => x"d4cdc287",
   196 => x"48d0ff58",
   197 => x"d4ff78c2",
   198 => x"78ffc348",
   199 => x"edf748c1",
   200 => x"5b5e0e87",
   201 => x"710e5d5c",
   202 => x"c54cc04b",
   203 => x"4adfcdee",
   204 => x"c348d4ff",
   205 => x"486878ff",
   206 => x"05a8fec3",
   207 => x"ff87fec0",
   208 => x"9b734dd4",
   209 => x"d087cc02",
   210 => x"49731e66",
   211 => x"c487e8f5",
   212 => x"ff87d686",
   213 => x"d1c448d0",
   214 => x"7dffc378",
   215 => x"c14866d0",
   216 => x"58a6d488",
   217 => x"f0059870",
   218 => x"48d4ff87",
   219 => x"7878ffc3",
   220 => x"c5059b73",
   221 => x"48d0ff87",
   222 => x"4ac178d0",
   223 => x"058ac14c",
   224 => x"7487edfe",
   225 => x"87c2f648",
   226 => x"711e731e",
   227 => x"ff4bc04a",
   228 => x"ffc348d4",
   229 => x"48d0ff78",
   230 => x"ff78c3c4",
   231 => x"ffc348d4",
   232 => x"c01e7278",
   233 => x"d1c1f0ff",
   234 => x"87e6f549",
   235 => x"987086c4",
   236 => x"c887d205",
   237 => x"66cc1ec0",
   238 => x"87e5fd49",
   239 => x"4b7086c4",
   240 => x"c248d0ff",
   241 => x"f5487378",
   242 => x"5e0e87c4",
   243 => x"0e5d5c5b",
   244 => x"ffc01ec0",
   245 => x"49c9c1f0",
   246 => x"d287f7f4",
   247 => x"d4cdc21e",
   248 => x"87fdfc49",
   249 => x"4cc086c8",
   250 => x"b7d284c1",
   251 => x"87f804ac",
   252 => x"97d4cdc2",
   253 => x"c0c349bf",
   254 => x"a9c0c199",
   255 => x"87e7c005",
   256 => x"97dbcdc2",
   257 => x"31d049bf",
   258 => x"97dccdc2",
   259 => x"32c84abf",
   260 => x"cdc2b172",
   261 => x"4abf97dd",
   262 => x"cf4c71b1",
   263 => x"9cffffff",
   264 => x"34ca84c1",
   265 => x"c287e7c1",
   266 => x"bf97ddcd",
   267 => x"c631c149",
   268 => x"decdc299",
   269 => x"c74abf97",
   270 => x"b1722ab7",
   271 => x"97d9cdc2",
   272 => x"cf4d4abf",
   273 => x"dacdc29d",
   274 => x"c34abf97",
   275 => x"c232ca9a",
   276 => x"bf97dbcd",
   277 => x"7333c24b",
   278 => x"dccdc2b2",
   279 => x"c34bbf97",
   280 => x"b7c69bc0",
   281 => x"c2b2732b",
   282 => x"7148c181",
   283 => x"c1497030",
   284 => x"70307548",
   285 => x"c14c724d",
   286 => x"c8947184",
   287 => x"06adb7c0",
   288 => x"34c187cc",
   289 => x"c0c82db7",
   290 => x"ff01adb7",
   291 => x"487487f4",
   292 => x"0e87f7f1",
   293 => x"5d5c5b5e",
   294 => x"c286f80e",
   295 => x"c048fad5",
   296 => x"f2cdc278",
   297 => x"fb49c01e",
   298 => x"86c487de",
   299 => x"c5059870",
   300 => x"c948c087",
   301 => x"4dc087c0",
   302 => x"edc07ec1",
   303 => x"c249bfe6",
   304 => x"714ae8ce",
   305 => x"e0ee4bc8",
   306 => x"05987087",
   307 => x"7ec087c2",
   308 => x"bfe2edc0",
   309 => x"c4cfc249",
   310 => x"4bc8714a",
   311 => x"7087caee",
   312 => x"87c20598",
   313 => x"026e7ec0",
   314 => x"c287fdc0",
   315 => x"4dbff8d4",
   316 => x"9ff0d5c2",
   317 => x"c5487ebf",
   318 => x"05a8ead6",
   319 => x"d4c287c7",
   320 => x"ce4dbff8",
   321 => x"ca486e87",
   322 => x"02a8d5e9",
   323 => x"48c087c5",
   324 => x"c287e3c7",
   325 => x"751ef2cd",
   326 => x"87ecf949",
   327 => x"987086c4",
   328 => x"c087c505",
   329 => x"87cec748",
   330 => x"bfe2edc0",
   331 => x"c4cfc249",
   332 => x"4bc8714a",
   333 => x"7087f2ec",
   334 => x"87c80598",
   335 => x"48fad5c2",
   336 => x"87da78c1",
   337 => x"bfe6edc0",
   338 => x"e8cec249",
   339 => x"4bc8714a",
   340 => x"7087d6ec",
   341 => x"c5c00298",
   342 => x"c648c087",
   343 => x"d5c287d8",
   344 => x"49bf97f0",
   345 => x"05a9d5c1",
   346 => x"c287cdc0",
   347 => x"bf97f1d5",
   348 => x"a9eac249",
   349 => x"87c5c002",
   350 => x"f9c548c0",
   351 => x"f2cdc287",
   352 => x"487ebf97",
   353 => x"02a8e9c3",
   354 => x"6e87cec0",
   355 => x"a8ebc348",
   356 => x"87c5c002",
   357 => x"ddc548c0",
   358 => x"fdcdc287",
   359 => x"9949bf97",
   360 => x"87ccc005",
   361 => x"97fecdc2",
   362 => x"a9c249bf",
   363 => x"87c5c002",
   364 => x"c1c548c0",
   365 => x"ffcdc287",
   366 => x"c248bf97",
   367 => x"7058f6d5",
   368 => x"88c1484c",
   369 => x"58fad5c2",
   370 => x"97c0cec2",
   371 => x"817549bf",
   372 => x"97c1cec2",
   373 => x"32c84abf",
   374 => x"c27ea172",
   375 => x"6e48c7da",
   376 => x"c2cec278",
   377 => x"c848bf97",
   378 => x"d5c258a6",
   379 => x"c202bffa",
   380 => x"edc087cf",
   381 => x"c249bfe2",
   382 => x"714ac4cf",
   383 => x"e8e94bc8",
   384 => x"02987087",
   385 => x"c087c5c0",
   386 => x"87eac348",
   387 => x"bff2d5c2",
   388 => x"dbdac24c",
   389 => x"d7cec25c",
   390 => x"c849bf97",
   391 => x"d6cec231",
   392 => x"a14abf97",
   393 => x"d8cec249",
   394 => x"d04abf97",
   395 => x"49a17232",
   396 => x"97d9cec2",
   397 => x"32d84abf",
   398 => x"c449a172",
   399 => x"dac29166",
   400 => x"c281bfc7",
   401 => x"c259cfda",
   402 => x"bf97dfce",
   403 => x"c232c84a",
   404 => x"bf97dece",
   405 => x"c24aa24b",
   406 => x"bf97e0ce",
   407 => x"7333d04b",
   408 => x"cec24aa2",
   409 => x"4bbf97e1",
   410 => x"33d89bcf",
   411 => x"c24aa273",
   412 => x"c25ad3da",
   413 => x"c292748a",
   414 => x"7248d3da",
   415 => x"c1c178a1",
   416 => x"c4cec287",
   417 => x"c849bf97",
   418 => x"c3cec231",
   419 => x"a14abf97",
   420 => x"c731c549",
   421 => x"29c981ff",
   422 => x"59dbdac2",
   423 => x"97c9cec2",
   424 => x"32c84abf",
   425 => x"97c8cec2",
   426 => x"4aa24bbf",
   427 => x"6e9266c4",
   428 => x"d7dac282",
   429 => x"cfdac25a",
   430 => x"c278c048",
   431 => x"7248cbda",
   432 => x"dac278a1",
   433 => x"dac248db",
   434 => x"c278bfcf",
   435 => x"c248dfda",
   436 => x"78bfd3da",
   437 => x"bffad5c2",
   438 => x"87c9c002",
   439 => x"30c44874",
   440 => x"c9c07e70",
   441 => x"d7dac287",
   442 => x"30c448bf",
   443 => x"d5c27e70",
   444 => x"786e48fe",
   445 => x"8ef848c1",
   446 => x"4c264d26",
   447 => x"4f264b26",
   448 => x"5c5b5e0e",
   449 => x"4a710e5d",
   450 => x"bffad5c2",
   451 => x"7287cb02",
   452 => x"722bc74b",
   453 => x"9dffc14d",
   454 => x"4b7287c9",
   455 => x"4d722bc8",
   456 => x"c29dffc3",
   457 => x"83bfc7da",
   458 => x"bfdeedc0",
   459 => x"87d902ab",
   460 => x"5be2edc0",
   461 => x"1ef2cdc2",
   462 => x"cbf14973",
   463 => x"7086c487",
   464 => x"87c50598",
   465 => x"e6c048c0",
   466 => x"fad5c287",
   467 => x"87d202bf",
   468 => x"91c44975",
   469 => x"81f2cdc2",
   470 => x"ffcf4c69",
   471 => x"9cffffff",
   472 => x"497587cb",
   473 => x"cdc291c2",
   474 => x"699f81f2",
   475 => x"fe48744c",
   476 => x"5e0e87c6",
   477 => x"0e5d5c5b",
   478 => x"4c7186f8",
   479 => x"87c5059c",
   480 => x"c0c348c0",
   481 => x"7ea4c887",
   482 => x"d878c048",
   483 => x"87c70266",
   484 => x"bf9766d8",
   485 => x"c087c505",
   486 => x"87e9c248",
   487 => x"49c11ec0",
   488 => x"87e3c749",
   489 => x"4d7086c4",
   490 => x"c2c1029d",
   491 => x"c2d6c287",
   492 => x"4966d84a",
   493 => x"7087d7e2",
   494 => x"f2c00298",
   495 => x"d84a7587",
   496 => x"4bcb4966",
   497 => x"7087fce2",
   498 => x"e2c00298",
   499 => x"751ec087",
   500 => x"87c7029d",
   501 => x"c048a6c8",
   502 => x"c887c578",
   503 => x"78c148a6",
   504 => x"c64966c8",
   505 => x"86c487e1",
   506 => x"059d4d70",
   507 => x"7587fefe",
   508 => x"cec1029d",
   509 => x"49a5dc87",
   510 => x"7869486e",
   511 => x"c449a5da",
   512 => x"a4c448a6",
   513 => x"48699f78",
   514 => x"780866c4",
   515 => x"bffad5c2",
   516 => x"d487d202",
   517 => x"699f49a5",
   518 => x"ffffc049",
   519 => x"d0487199",
   520 => x"c27e7030",
   521 => x"6e7ec087",
   522 => x"bf66c448",
   523 => x"0866c480",
   524 => x"cc7cc078",
   525 => x"66c449a4",
   526 => x"a4d079bf",
   527 => x"c179c049",
   528 => x"c087c248",
   529 => x"fa8ef848",
   530 => x"5e0e87ee",
   531 => x"710e5c5b",
   532 => x"c1029c4c",
   533 => x"a4c887cb",
   534 => x"c1026949",
   535 => x"496c87c3",
   536 => x"714866cc",
   537 => x"58a6d080",
   538 => x"d5c2b970",
   539 => x"ff4abff6",
   540 => x"719972ba",
   541 => x"e5c00299",
   542 => x"4ba4c487",
   543 => x"fff9496b",
   544 => x"c27b7087",
   545 => x"49bff2d5",
   546 => x"7c71816c",
   547 => x"c2b966cc",
   548 => x"4abff6d5",
   549 => x"9972baff",
   550 => x"ff059971",
   551 => x"66cc87db",
   552 => x"87d6f97c",
   553 => x"711e731e",
   554 => x"c7029b4b",
   555 => x"49a3c887",
   556 => x"87c50569",
   557 => x"f6c048c0",
   558 => x"cbdac287",
   559 => x"a3c449bf",
   560 => x"c24a6a4a",
   561 => x"f2d5c28a",
   562 => x"a17292bf",
   563 => x"f6d5c249",
   564 => x"9a6b4abf",
   565 => x"c049a172",
   566 => x"c859e2ed",
   567 => x"ea711e66",
   568 => x"86c487e6",
   569 => x"c4059870",
   570 => x"c248c087",
   571 => x"f848c187",
   572 => x"731e87ca",
   573 => x"9b4b711e",
   574 => x"87e4c002",
   575 => x"5bdfdac2",
   576 => x"8ac24a73",
   577 => x"bff2d5c2",
   578 => x"dac29249",
   579 => x"7248bfcb",
   580 => x"e3dac280",
   581 => x"c4487158",
   582 => x"c2d6c230",
   583 => x"87edc058",
   584 => x"48dbdac2",
   585 => x"bfcfdac2",
   586 => x"dfdac278",
   587 => x"d3dac248",
   588 => x"d5c278bf",
   589 => x"c902bffa",
   590 => x"f2d5c287",
   591 => x"31c449bf",
   592 => x"dac287c7",
   593 => x"c449bfd7",
   594 => x"c2d6c231",
   595 => x"87ecf659",
   596 => x"5c5b5e0e",
   597 => x"c04a710e",
   598 => x"029a724b",
   599 => x"da87e0c0",
   600 => x"699f49a2",
   601 => x"fad5c24b",
   602 => x"87cf02bf",
   603 => x"9f49a2d4",
   604 => x"c04c4969",
   605 => x"d09cffff",
   606 => x"c087c234",
   607 => x"73b3744c",
   608 => x"87eefd49",
   609 => x"0e87f3f5",
   610 => x"5d5c5b5e",
   611 => x"7186f40e",
   612 => x"727ec04a",
   613 => x"87d8029a",
   614 => x"48eecdc2",
   615 => x"cdc278c0",
   616 => x"dac248e6",
   617 => x"c278bfdf",
   618 => x"c248eacd",
   619 => x"78bfdbda",
   620 => x"48cfd6c2",
   621 => x"d5c250c0",
   622 => x"c249bffe",
   623 => x"4abfeecd",
   624 => x"c403aa71",
   625 => x"497287c9",
   626 => x"c00599cf",
   627 => x"edc087e9",
   628 => x"cdc248de",
   629 => x"c278bfe6",
   630 => x"c21ef2cd",
   631 => x"49bfe6cd",
   632 => x"48e6cdc2",
   633 => x"7178a1c1",
   634 => x"c487dde6",
   635 => x"daedc086",
   636 => x"f2cdc248",
   637 => x"c087cc78",
   638 => x"48bfdaed",
   639 => x"c080e0c0",
   640 => x"c258deed",
   641 => x"48bfeecd",
   642 => x"cdc280c1",
   643 => x"5a2758f2",
   644 => x"bf00000b",
   645 => x"9d4dbf97",
   646 => x"87e3c202",
   647 => x"02ade5c3",
   648 => x"c087dcc2",
   649 => x"4bbfdaed",
   650 => x"1149a3cb",
   651 => x"05accf4c",
   652 => x"7587d2c1",
   653 => x"c199df49",
   654 => x"c291cd89",
   655 => x"c181c2d6",
   656 => x"51124aa3",
   657 => x"124aa3c3",
   658 => x"4aa3c551",
   659 => x"a3c75112",
   660 => x"c951124a",
   661 => x"51124aa3",
   662 => x"124aa3ce",
   663 => x"4aa3d051",
   664 => x"a3d25112",
   665 => x"d451124a",
   666 => x"51124aa3",
   667 => x"124aa3d6",
   668 => x"4aa3d851",
   669 => x"a3dc5112",
   670 => x"de51124a",
   671 => x"51124aa3",
   672 => x"fac07ec1",
   673 => x"c8497487",
   674 => x"ebc00599",
   675 => x"d0497487",
   676 => x"87d10599",
   677 => x"c00266dc",
   678 => x"497387cb",
   679 => x"700f66dc",
   680 => x"d3c00298",
   681 => x"c0056e87",
   682 => x"d6c287c6",
   683 => x"50c048c2",
   684 => x"bfdaedc0",
   685 => x"87ddc248",
   686 => x"48cfd6c2",
   687 => x"c27e50c0",
   688 => x"49bffed5",
   689 => x"bfeecdc2",
   690 => x"04aa714a",
   691 => x"c287f7fb",
   692 => x"05bfdfda",
   693 => x"c287c8c0",
   694 => x"02bffad5",
   695 => x"c287f4c1",
   696 => x"49bfeacd",
   697 => x"c287d9f0",
   698 => x"c458eecd",
   699 => x"cdc248a6",
   700 => x"c278bfea",
   701 => x"02bffad5",
   702 => x"c487d8c0",
   703 => x"ffcf4966",
   704 => x"99f8ffff",
   705 => x"c5c002a9",
   706 => x"c04cc087",
   707 => x"4cc187e1",
   708 => x"c487dcc0",
   709 => x"ffcf4966",
   710 => x"02a999f8",
   711 => x"c887c8c0",
   712 => x"78c048a6",
   713 => x"c887c5c0",
   714 => x"78c148a6",
   715 => x"744c66c8",
   716 => x"dec0059c",
   717 => x"4966c487",
   718 => x"d5c289c2",
   719 => x"c291bff2",
   720 => x"48bfcbda",
   721 => x"cdc28071",
   722 => x"cdc258ea",
   723 => x"78c048ee",
   724 => x"c087e3f9",
   725 => x"ee8ef448",
   726 => x"000087de",
   727 => x"ffff0000",
   728 => x"0b6affff",
   729 => x"0b730000",
   730 => x"41460000",
   731 => x"20323354",
   732 => x"46002020",
   733 => x"36315441",
   734 => x"00202020",
   735 => x"48d4ff1e",
   736 => x"6878ffc3",
   737 => x"1e4f2648",
   738 => x"c348d4ff",
   739 => x"d0ff78ff",
   740 => x"78e1c048",
   741 => x"d448d4ff",
   742 => x"e3dac278",
   743 => x"bfd4ff48",
   744 => x"1e4f2650",
   745 => x"c048d0ff",
   746 => x"4f2678e0",
   747 => x"87ccff1e",
   748 => x"02994970",
   749 => x"fbc087c6",
   750 => x"87f105a9",
   751 => x"4f264871",
   752 => x"5c5b5e0e",
   753 => x"c04b710e",
   754 => x"87f0fe4c",
   755 => x"02994970",
   756 => x"c087f9c0",
   757 => x"c002a9ec",
   758 => x"fbc087f2",
   759 => x"ebc002a9",
   760 => x"b766cc87",
   761 => x"87c703ac",
   762 => x"c20266d0",
   763 => x"71537187",
   764 => x"87c20299",
   765 => x"c3fe84c1",
   766 => x"99497087",
   767 => x"c087cd02",
   768 => x"c702a9ec",
   769 => x"a9fbc087",
   770 => x"87d5ff05",
   771 => x"c30266d0",
   772 => x"7b97c087",
   773 => x"05a9ecc0",
   774 => x"4a7487c4",
   775 => x"4a7487c5",
   776 => x"728a0ac0",
   777 => x"2687c248",
   778 => x"264c264d",
   779 => x"1e4f264b",
   780 => x"7087c9fd",
   781 => x"aaf0c04a",
   782 => x"c087c904",
   783 => x"c301aaf9",
   784 => x"8af0c087",
   785 => x"04aac1c1",
   786 => x"dac187c9",
   787 => x"87c301aa",
   788 => x"728af7c0",
   789 => x"0e4f2648",
   790 => x"0e5c5b5e",
   791 => x"d4ff4a71",
   792 => x"c049724b",
   793 => x"4c7087e7",
   794 => x"87c2029c",
   795 => x"d0ff8cc1",
   796 => x"c178c548",
   797 => x"49747bd5",
   798 => x"dec131c6",
   799 => x"4abf97c0",
   800 => x"70b07148",
   801 => x"48d0ff7b",
   802 => x"dcfe78c4",
   803 => x"5b5e0e87",
   804 => x"f80e5d5c",
   805 => x"c04c7186",
   806 => x"87ebfb7e",
   807 => x"f4c04bc0",
   808 => x"49bf97fa",
   809 => x"cf04a9c0",
   810 => x"87c0fc87",
   811 => x"f4c083c1",
   812 => x"49bf97fa",
   813 => x"87f106ab",
   814 => x"97faf4c0",
   815 => x"87cf02bf",
   816 => x"7087f9fa",
   817 => x"c6029949",
   818 => x"a9ecc087",
   819 => x"c087f105",
   820 => x"87e8fa4b",
   821 => x"e3fa4d70",
   822 => x"58a6c887",
   823 => x"7087ddfa",
   824 => x"c883c14a",
   825 => x"699749a4",
   826 => x"c702ad49",
   827 => x"adffc087",
   828 => x"87e7c005",
   829 => x"9749a4c9",
   830 => x"66c44969",
   831 => x"87c702a9",
   832 => x"a8ffc048",
   833 => x"ca87d405",
   834 => x"699749a4",
   835 => x"c602aa49",
   836 => x"aaffc087",
   837 => x"c187c405",
   838 => x"c087d07e",
   839 => x"c602adec",
   840 => x"adfbc087",
   841 => x"c087c405",
   842 => x"6e7ec14b",
   843 => x"87e1fe02",
   844 => x"7387f0f9",
   845 => x"fb8ef848",
   846 => x"0e0087ed",
   847 => x"5d5c5b5e",
   848 => x"7186f80e",
   849 => x"4bd4ff4d",
   850 => x"dac21e75",
   851 => x"e1e849e8",
   852 => x"7086c487",
   853 => x"cac40298",
   854 => x"48a6c487",
   855 => x"bfc2dec1",
   856 => x"fb497578",
   857 => x"d0ff87f1",
   858 => x"c178c548",
   859 => x"4ac07bd6",
   860 => x"1149a275",
   861 => x"cb82c17b",
   862 => x"f304aab7",
   863 => x"c34acc87",
   864 => x"82c17bff",
   865 => x"aab7e0c0",
   866 => x"ff87f404",
   867 => x"78c448d0",
   868 => x"c57bffc3",
   869 => x"7bd3c178",
   870 => x"78c47bc1",
   871 => x"b7c04866",
   872 => x"eec206a8",
   873 => x"f0dac287",
   874 => x"66c44cbf",
   875 => x"c8887448",
   876 => x"9c7458a6",
   877 => x"87f7c102",
   878 => x"7ef2cdc2",
   879 => x"8c4dc0c8",
   880 => x"03acb7c0",
   881 => x"c0c887c6",
   882 => x"4cc04da4",
   883 => x"97e3dac2",
   884 => x"99d049bf",
   885 => x"c087d002",
   886 => x"e8dac21e",
   887 => x"87c4eb49",
   888 => x"4a7086c4",
   889 => x"c287edc0",
   890 => x"c21ef2cd",
   891 => x"ea49e8da",
   892 => x"86c487f2",
   893 => x"d0ff4a70",
   894 => x"78c5c848",
   895 => x"6e7bd4c1",
   896 => x"6e7bbf97",
   897 => x"7080c148",
   898 => x"058dc17e",
   899 => x"ff87f0ff",
   900 => x"78c448d0",
   901 => x"c5059a72",
   902 => x"c148c087",
   903 => x"1ec187c7",
   904 => x"49e8dac2",
   905 => x"c487e3e8",
   906 => x"059c7486",
   907 => x"c487c9fe",
   908 => x"b7c04866",
   909 => x"87d106a8",
   910 => x"48e8dac2",
   911 => x"80d078c0",
   912 => x"80f478c0",
   913 => x"bff4dac2",
   914 => x"4866c478",
   915 => x"01a8b7c0",
   916 => x"ff87d2fd",
   917 => x"78c548d0",
   918 => x"c07bd3c1",
   919 => x"c178c47b",
   920 => x"c087c248",
   921 => x"268ef848",
   922 => x"264c264d",
   923 => x"0e4f264b",
   924 => x"5d5c5b5e",
   925 => x"4b711e0e",
   926 => x"ab4d4cc0",
   927 => x"87e8c004",
   928 => x"1ecdf2c0",
   929 => x"c4029d75",
   930 => x"c24ac087",
   931 => x"724ac187",
   932 => x"87f3eb49",
   933 => x"7e7086c4",
   934 => x"056e84c1",
   935 => x"4c7387c2",
   936 => x"ac7385c1",
   937 => x"87d8ff06",
   938 => x"fe26486e",
   939 => x"711e87f9",
   940 => x"0566c44a",
   941 => x"497287c5",
   942 => x"2687c0fa",
   943 => x"5b5e0e4f",
   944 => x"1e0e5d5c",
   945 => x"de494c71",
   946 => x"d0dbc291",
   947 => x"9785714d",
   948 => x"dcc1026d",
   949 => x"fcdac287",
   950 => x"817449bf",
   951 => x"87cffe71",
   952 => x"98487e70",
   953 => x"87f2c002",
   954 => x"4bc4dbc2",
   955 => x"49cb4a70",
   956 => x"87f3c6ff",
   957 => x"93cb4b74",
   958 => x"83d4dec1",
   959 => x"fcc083c4",
   960 => x"49747bf5",
   961 => x"87f6c0c1",
   962 => x"dec17b75",
   963 => x"49bf97c1",
   964 => x"c4dbc21e",
   965 => x"87d6fe49",
   966 => x"497486c4",
   967 => x"87dec0c1",
   968 => x"c1c149c0",
   969 => x"dac287fd",
   970 => x"78c048e4",
   971 => x"f9dd49c1",
   972 => x"f2fc2687",
   973 => x"616f4c87",
   974 => x"676e6964",
   975 => x"002e2e2e",
   976 => x"711e731e",
   977 => x"dac2494a",
   978 => x"7181bffc",
   979 => x"7087e0fc",
   980 => x"c4029b4b",
   981 => x"f7e74987",
   982 => x"fcdac287",
   983 => x"c178c048",
   984 => x"87c6dd49",
   985 => x"1e87c4fc",
   986 => x"c0c149c0",
   987 => x"4f2687f5",
   988 => x"494a711e",
   989 => x"dec191cb",
   990 => x"81c881d4",
   991 => x"dac24811",
   992 => x"dac258e8",
   993 => x"78c048fc",
   994 => x"dddc49c1",
   995 => x"1e4f2687",
   996 => x"d2029971",
   997 => x"e9dfc187",
   998 => x"f750c048",
   999 => x"f0fdc080",
  1000 => x"cddec140",
  1001 => x"c187ce78",
  1002 => x"c148e5df",
  1003 => x"fc78c6de",
  1004 => x"e7fdc080",
  1005 => x"0e4f2678",
  1006 => x"5d5c5b5e",
  1007 => x"c286f40e",
  1008 => x"c04df2cd",
  1009 => x"48a6c44c",
  1010 => x"dac278c0",
  1011 => x"c048bffc",
  1012 => x"c0c106a8",
  1013 => x"f2cdc287",
  1014 => x"c0029848",
  1015 => x"f2c087f7",
  1016 => x"66c81ecd",
  1017 => x"c487c702",
  1018 => x"78c048a6",
  1019 => x"a6c487c5",
  1020 => x"c478c148",
  1021 => x"cee64966",
  1022 => x"7086c487",
  1023 => x"c484c14d",
  1024 => x"80c14866",
  1025 => x"c258a6c8",
  1026 => x"acbffcda",
  1027 => x"7587c603",
  1028 => x"c9ff059d",
  1029 => x"754cc087",
  1030 => x"dcc3029d",
  1031 => x"cdf2c087",
  1032 => x"0266c81e",
  1033 => x"a6cc87c7",
  1034 => x"c578c048",
  1035 => x"48a6cc87",
  1036 => x"66cc78c1",
  1037 => x"87cfe549",
  1038 => x"7e7086c4",
  1039 => x"c2029848",
  1040 => x"cb4987e4",
  1041 => x"49699781",
  1042 => x"c10299d0",
  1043 => x"497487d4",
  1044 => x"dec191cb",
  1045 => x"fdc081d4",
  1046 => x"81c879c0",
  1047 => x"7451ffc3",
  1048 => x"c291de49",
  1049 => x"714dd0db",
  1050 => x"97c1c285",
  1051 => x"49a5c17d",
  1052 => x"c251e0c0",
  1053 => x"bf97c2d6",
  1054 => x"c187d202",
  1055 => x"4ba5c284",
  1056 => x"4ac2d6c2",
  1057 => x"c0ff49db",
  1058 => x"d9c187dd",
  1059 => x"49a5cd87",
  1060 => x"84c151c0",
  1061 => x"6e4ba5c2",
  1062 => x"ff49cb4a",
  1063 => x"c187c8c0",
  1064 => x"497487c4",
  1065 => x"dec191cb",
  1066 => x"fac081d4",
  1067 => x"d6c279fd",
  1068 => x"02bf97c2",
  1069 => x"497487d8",
  1070 => x"84c191de",
  1071 => x"4bd0dbc2",
  1072 => x"d6c28371",
  1073 => x"49dd4ac2",
  1074 => x"87dbfffe",
  1075 => x"4b7487d8",
  1076 => x"dbc293de",
  1077 => x"a3cb83d0",
  1078 => x"c151c049",
  1079 => x"4a6e7384",
  1080 => x"fffe49cb",
  1081 => x"66c487c1",
  1082 => x"c880c148",
  1083 => x"acc758a6",
  1084 => x"87c5c003",
  1085 => x"e4fc056e",
  1086 => x"f4487487",
  1087 => x"87e7f58e",
  1088 => x"711e731e",
  1089 => x"91cb494b",
  1090 => x"81d4dec1",
  1091 => x"c14aa1c8",
  1092 => x"1248c0de",
  1093 => x"4aa1c950",
  1094 => x"48faf4c0",
  1095 => x"81ca5012",
  1096 => x"48c1dec1",
  1097 => x"dec15011",
  1098 => x"49bf97c1",
  1099 => x"f549c01e",
  1100 => x"dac287fc",
  1101 => x"78de48e4",
  1102 => x"edd549c1",
  1103 => x"eaf42687",
  1104 => x"5b5e0e87",
  1105 => x"f40e5d5c",
  1106 => x"494d7186",
  1107 => x"dec191cb",
  1108 => x"a1c881d4",
  1109 => x"7ea1ca4a",
  1110 => x"c248a6c4",
  1111 => x"78bfecde",
  1112 => x"4bbf976e",
  1113 => x"734c66c4",
  1114 => x"cc48122c",
  1115 => x"9c7058a6",
  1116 => x"81c984c1",
  1117 => x"b7496997",
  1118 => x"87c204ac",
  1119 => x"976e4cc0",
  1120 => x"66c84abf",
  1121 => x"ff317249",
  1122 => x"9966c4b9",
  1123 => x"30724874",
  1124 => x"71484a70",
  1125 => x"f0dec2b0",
  1126 => x"e1e4c058",
  1127 => x"d449c087",
  1128 => x"497587c8",
  1129 => x"87d6f6c0",
  1130 => x"faf28ef4",
  1131 => x"1e731e87",
  1132 => x"fe494b71",
  1133 => x"497387cb",
  1134 => x"f287c6fe",
  1135 => x"731e87ed",
  1136 => x"c64b711e",
  1137 => x"db024aa3",
  1138 => x"028ac187",
  1139 => x"028a87d6",
  1140 => x"8a87dac1",
  1141 => x"87fcc002",
  1142 => x"e1c0028a",
  1143 => x"cb028a87",
  1144 => x"87dbc187",
  1145 => x"c7f649c7",
  1146 => x"87dec187",
  1147 => x"bffcdac2",
  1148 => x"87cbc102",
  1149 => x"c288c148",
  1150 => x"c158c0db",
  1151 => x"dbc287c1",
  1152 => x"c002bfc0",
  1153 => x"dac287f9",
  1154 => x"c148bffc",
  1155 => x"c0dbc280",
  1156 => x"87ebc058",
  1157 => x"bffcdac2",
  1158 => x"c289c649",
  1159 => x"c059c0db",
  1160 => x"da03a9b7",
  1161 => x"fcdac287",
  1162 => x"d278c048",
  1163 => x"c0dbc287",
  1164 => x"87cb02bf",
  1165 => x"bffcdac2",
  1166 => x"c280c648",
  1167 => x"c058c0db",
  1168 => x"87e6d149",
  1169 => x"f3c04973",
  1170 => x"def087f4",
  1171 => x"5b5e0e87",
  1172 => x"ff0e5d5c",
  1173 => x"a6dc86d4",
  1174 => x"48a6c859",
  1175 => x"80c478c0",
  1176 => x"7866c0c1",
  1177 => x"78c180c4",
  1178 => x"78c180c4",
  1179 => x"48c0dbc2",
  1180 => x"dac278c1",
  1181 => x"de48bfe4",
  1182 => x"87c905a8",
  1183 => x"cc87f8f4",
  1184 => x"e4cf58a6",
  1185 => x"87ffe387",
  1186 => x"e387e1e4",
  1187 => x"4c7087ee",
  1188 => x"02acfbc0",
  1189 => x"d887fbc1",
  1190 => x"edc10566",
  1191 => x"66fcc087",
  1192 => x"6a82c44a",
  1193 => x"c11e727e",
  1194 => x"c448deda",
  1195 => x"a1c84966",
  1196 => x"7141204a",
  1197 => x"87f905aa",
  1198 => x"4a265110",
  1199 => x"4866fcc0",
  1200 => x"78c0c4c1",
  1201 => x"81c7496a",
  1202 => x"fcc05174",
  1203 => x"81c84966",
  1204 => x"fcc051c1",
  1205 => x"81c94966",
  1206 => x"fcc051c0",
  1207 => x"81ca4966",
  1208 => x"1ec151c0",
  1209 => x"496a1ed8",
  1210 => x"d3e381c8",
  1211 => x"c186c887",
  1212 => x"c04866c0",
  1213 => x"87c701a8",
  1214 => x"c148a6c8",
  1215 => x"c187ce78",
  1216 => x"c14866c0",
  1217 => x"58a6d088",
  1218 => x"dfe287c3",
  1219 => x"48a6d087",
  1220 => x"9c7478c2",
  1221 => x"87cdcd02",
  1222 => x"c14866c8",
  1223 => x"03a866c4",
  1224 => x"dc87c2cd",
  1225 => x"78c048a6",
  1226 => x"78c080e8",
  1227 => x"7087cde1",
  1228 => x"acd0c14c",
  1229 => x"87d5c205",
  1230 => x"e37e66c4",
  1231 => x"a6c887f1",
  1232 => x"87f8e058",
  1233 => x"ecc04c70",
  1234 => x"ebc105ac",
  1235 => x"4966c887",
  1236 => x"fcc091cb",
  1237 => x"a1c48166",
  1238 => x"c84d6a4a",
  1239 => x"66c44aa1",
  1240 => x"f0fdc052",
  1241 => x"87d4e079",
  1242 => x"029c4c70",
  1243 => x"fbc087d8",
  1244 => x"87d202ac",
  1245 => x"c3e05574",
  1246 => x"9c4c7087",
  1247 => x"c087c702",
  1248 => x"ff05acfb",
  1249 => x"e0c087ee",
  1250 => x"55c1c255",
  1251 => x"d87d97c0",
  1252 => x"a86e4866",
  1253 => x"c887db05",
  1254 => x"66cc4866",
  1255 => x"87ca04a8",
  1256 => x"c14866c8",
  1257 => x"58a6cc80",
  1258 => x"66cc87c8",
  1259 => x"d088c148",
  1260 => x"dfff58a6",
  1261 => x"4c7087c6",
  1262 => x"05acd0c1",
  1263 => x"66d487c8",
  1264 => x"d880c148",
  1265 => x"d0c158a6",
  1266 => x"ebfd02ac",
  1267 => x"4866c487",
  1268 => x"05a866d8",
  1269 => x"c087e0c9",
  1270 => x"c048a6e0",
  1271 => x"c0487478",
  1272 => x"7e7088fb",
  1273 => x"c9029848",
  1274 => x"cb4887e2",
  1275 => x"487e7088",
  1276 => x"cdc10298",
  1277 => x"88c94887",
  1278 => x"98487e70",
  1279 => x"87fec302",
  1280 => x"7088c448",
  1281 => x"0298487e",
  1282 => x"c14887ce",
  1283 => x"487e7088",
  1284 => x"e9c30298",
  1285 => x"87d6c887",
  1286 => x"c048a6dc",
  1287 => x"ddff78f0",
  1288 => x"4c7087da",
  1289 => x"02acecc0",
  1290 => x"c087c4c0",
  1291 => x"c05ca6e0",
  1292 => x"cd02acec",
  1293 => x"c3ddff87",
  1294 => x"c04c7087",
  1295 => x"ff05acec",
  1296 => x"ecc087f3",
  1297 => x"c4c002ac",
  1298 => x"efdcff87",
  1299 => x"ca1ec087",
  1300 => x"4966d01e",
  1301 => x"c4c191cb",
  1302 => x"80714866",
  1303 => x"c858a6cc",
  1304 => x"80c44866",
  1305 => x"cc58a6d0",
  1306 => x"ff49bf66",
  1307 => x"c187d1dd",
  1308 => x"d41ede1e",
  1309 => x"ff49bf66",
  1310 => x"d087c5dd",
  1311 => x"48497086",
  1312 => x"c08808c0",
  1313 => x"c058a6e8",
  1314 => x"eec006a8",
  1315 => x"66e4c087",
  1316 => x"03a8dd48",
  1317 => x"c487e4c0",
  1318 => x"c049bf66",
  1319 => x"c08166e4",
  1320 => x"e4c051e0",
  1321 => x"81c14966",
  1322 => x"81bf66c4",
  1323 => x"c051c1c2",
  1324 => x"c24966e4",
  1325 => x"bf66c481",
  1326 => x"6e51c081",
  1327 => x"c0c4c148",
  1328 => x"c8496e78",
  1329 => x"5166d081",
  1330 => x"81c9496e",
  1331 => x"6e5166d4",
  1332 => x"dc81ca49",
  1333 => x"66d05166",
  1334 => x"d480c148",
  1335 => x"66c858a6",
  1336 => x"a866cc48",
  1337 => x"87cbc004",
  1338 => x"c14866c8",
  1339 => x"58a6cc80",
  1340 => x"cc87d9c5",
  1341 => x"88c14866",
  1342 => x"c558a6d0",
  1343 => x"dcff87ce",
  1344 => x"e8c087ed",
  1345 => x"dcff58a6",
  1346 => x"e0c087e5",
  1347 => x"ecc058a6",
  1348 => x"cac005a8",
  1349 => x"48a6dc87",
  1350 => x"7866e4c0",
  1351 => x"ff87c4c0",
  1352 => x"c887d9d9",
  1353 => x"91cb4966",
  1354 => x"4866fcc0",
  1355 => x"7e708071",
  1356 => x"6e82c84a",
  1357 => x"c081ca49",
  1358 => x"dc5166e4",
  1359 => x"81c14966",
  1360 => x"8966e4c0",
  1361 => x"307148c1",
  1362 => x"89c14970",
  1363 => x"c27a9771",
  1364 => x"49bfecde",
  1365 => x"2966e4c0",
  1366 => x"484a6a97",
  1367 => x"ecc09871",
  1368 => x"496e58a6",
  1369 => x"4d6981c4",
  1370 => x"c44866d8",
  1371 => x"c002a866",
  1372 => x"a6c487c8",
  1373 => x"c078c048",
  1374 => x"a6c487c5",
  1375 => x"c478c148",
  1376 => x"e0c01e66",
  1377 => x"ff49751e",
  1378 => x"c887f5d8",
  1379 => x"c04c7086",
  1380 => x"c106acb7",
  1381 => x"857487d4",
  1382 => x"7449e0c0",
  1383 => x"c14b7589",
  1384 => x"714ae7da",
  1385 => x"87ffebfe",
  1386 => x"e0c085c2",
  1387 => x"80c14866",
  1388 => x"58a6e4c0",
  1389 => x"4966e8c0",
  1390 => x"a97081c1",
  1391 => x"87c8c002",
  1392 => x"c048a6c4",
  1393 => x"87c5c078",
  1394 => x"c148a6c4",
  1395 => x"1e66c478",
  1396 => x"c049a4c2",
  1397 => x"887148e0",
  1398 => x"751e4970",
  1399 => x"dfd7ff49",
  1400 => x"c086c887",
  1401 => x"ff01a8b7",
  1402 => x"e0c087c0",
  1403 => x"d1c00266",
  1404 => x"c9496e87",
  1405 => x"66e0c081",
  1406 => x"c1486e51",
  1407 => x"c078c1c5",
  1408 => x"496e87cc",
  1409 => x"51c281c9",
  1410 => x"c6c1486e",
  1411 => x"66c878ed",
  1412 => x"a866cc48",
  1413 => x"87cbc004",
  1414 => x"c14866c8",
  1415 => x"58a6cc80",
  1416 => x"cc87e9c0",
  1417 => x"88c14866",
  1418 => x"c058a6d0",
  1419 => x"d5ff87de",
  1420 => x"4c7087fa",
  1421 => x"c187d5c0",
  1422 => x"c005acc6",
  1423 => x"66d087c8",
  1424 => x"d480c148",
  1425 => x"d5ff58a6",
  1426 => x"4c7087e2",
  1427 => x"c14866d4",
  1428 => x"58a6d880",
  1429 => x"c0029c74",
  1430 => x"66c887cb",
  1431 => x"66c4c148",
  1432 => x"fef204a8",
  1433 => x"fad4ff87",
  1434 => x"4866c887",
  1435 => x"c003a8c7",
  1436 => x"dbc287e5",
  1437 => x"78c048c0",
  1438 => x"cb4966c8",
  1439 => x"66fcc091",
  1440 => x"4aa1c481",
  1441 => x"52c04a6a",
  1442 => x"4866c879",
  1443 => x"a6cc80c1",
  1444 => x"04a8c758",
  1445 => x"ff87dbff",
  1446 => x"dfff8ed4",
  1447 => x"6f4c87c9",
  1448 => x"2a206461",
  1449 => x"3a00202e",
  1450 => x"731e0020",
  1451 => x"9b4b711e",
  1452 => x"c287c602",
  1453 => x"c048fcda",
  1454 => x"c21ec778",
  1455 => x"1ebffcda",
  1456 => x"1ed4dec1",
  1457 => x"bfe4dac2",
  1458 => x"87c1ee49",
  1459 => x"dac286cc",
  1460 => x"e249bfe4",
  1461 => x"9b7387f9",
  1462 => x"c187c802",
  1463 => x"c049d4de",
  1464 => x"ff87ede2",
  1465 => x"1e87c4de",
  1466 => x"48c0dec1",
  1467 => x"dfc150c0",
  1468 => x"ff49bff7",
  1469 => x"c087c4d9",
  1470 => x"1e4f2648",
  1471 => x"c187dfc7",
  1472 => x"87e6fe49",
  1473 => x"87e8eefe",
  1474 => x"cd029870",
  1475 => x"c2f6fe87",
  1476 => x"02987087",
  1477 => x"4ac187c4",
  1478 => x"4ac087c2",
  1479 => x"ce059a72",
  1480 => x"c11ec087",
  1481 => x"c049cbdd",
  1482 => x"c487dbee",
  1483 => x"c087fe86",
  1484 => x"d6ddc11e",
  1485 => x"cdeec049",
  1486 => x"fe1ec087",
  1487 => x"497087e9",
  1488 => x"87c2eec0",
  1489 => x"f887d6c3",
  1490 => x"534f268e",
  1491 => x"61662044",
  1492 => x"64656c69",
  1493 => x"6f42002e",
  1494 => x"6e69746f",
  1495 => x"2e2e2e67",
  1496 => x"e5c01e00",
  1497 => x"87fa87e7",
  1498 => x"c21e4f26",
  1499 => x"c048fcda",
  1500 => x"e4dac278",
  1501 => x"fe78c048",
  1502 => x"87e587c1",
  1503 => x"4f2648c0",
  1504 => x"00010000",
  1505 => x"20800000",
  1506 => x"74697845",
  1507 => x"42208000",
  1508 => x"006b6361",
  1509 => x"00000ebd",
  1510 => x"000026d0",
  1511 => x"bd000000",
  1512 => x"ee00000e",
  1513 => x"00000026",
  1514 => x"0ebd0000",
  1515 => x"270c0000",
  1516 => x"00000000",
  1517 => x"000ebd00",
  1518 => x"00272a00",
  1519 => x"00000000",
  1520 => x"00000ebd",
  1521 => x"00002748",
  1522 => x"bd000000",
  1523 => x"6600000e",
  1524 => x"00000027",
  1525 => x"0ebd0000",
  1526 => x"27840000",
  1527 => x"00000000",
  1528 => x"000f7000",
  1529 => x"00000000",
  1530 => x"00000000",
  1531 => x"000011be",
  1532 => x"00000000",
  1533 => x"fb000000",
  1534 => x"42000017",
  1535 => x"20544f4f",
  1536 => x"52202020",
  1537 => x"1e004d4f",
  1538 => x"c048f0fe",
  1539 => x"7909cd78",
  1540 => x"1e4f2609",
  1541 => x"bff0fe1e",
  1542 => x"2626487e",
  1543 => x"f0fe1e4f",
  1544 => x"2678c148",
  1545 => x"f0fe1e4f",
  1546 => x"2678c048",
  1547 => x"4a711e4f",
  1548 => x"265252c0",
  1549 => x"5b5e0e4f",
  1550 => x"f40e5d5c",
  1551 => x"974d7186",
  1552 => x"a5c17e6d",
  1553 => x"486c974c",
  1554 => x"6e58a6c8",
  1555 => x"a866c448",
  1556 => x"ff87c505",
  1557 => x"87e6c048",
  1558 => x"c287caff",
  1559 => x"6c9749a5",
  1560 => x"4ba3714b",
  1561 => x"974b6b97",
  1562 => x"486e7e6c",
  1563 => x"a6c880c1",
  1564 => x"cc98c758",
  1565 => x"977058a6",
  1566 => x"87e1fe7c",
  1567 => x"8ef44873",
  1568 => x"4c264d26",
  1569 => x"4f264b26",
  1570 => x"5c5b5e0e",
  1571 => x"7186f40e",
  1572 => x"4a66d84c",
  1573 => x"c29affc3",
  1574 => x"6c974ba4",
  1575 => x"49a17349",
  1576 => x"6c975172",
  1577 => x"c1486e7e",
  1578 => x"58a6c880",
  1579 => x"a6cc98c7",
  1580 => x"f4547058",
  1581 => x"87caff8e",
  1582 => x"e8fd1e1e",
  1583 => x"4abfe087",
  1584 => x"c0e0c049",
  1585 => x"87cb0299",
  1586 => x"dec21e72",
  1587 => x"f7fe49e2",
  1588 => x"fc86c487",
  1589 => x"7e7087fd",
  1590 => x"2687c2fd",
  1591 => x"c21e4f26",
  1592 => x"fd49e2de",
  1593 => x"e2c187c7",
  1594 => x"dafc49f8",
  1595 => x"87f7c387",
  1596 => x"5e0e4f26",
  1597 => x"0e5d5c5b",
  1598 => x"dec24d71",
  1599 => x"f4fc49e2",
  1600 => x"c04b7087",
  1601 => x"c304abb7",
  1602 => x"f0c387c2",
  1603 => x"87c905ab",
  1604 => x"48d6e7c1",
  1605 => x"e3c278c1",
  1606 => x"abe0c387",
  1607 => x"c187c905",
  1608 => x"c148dae7",
  1609 => x"87d4c278",
  1610 => x"bfdae7c1",
  1611 => x"c287c602",
  1612 => x"c24ca3c0",
  1613 => x"c14c7387",
  1614 => x"02bfd6e7",
  1615 => x"7487e0c0",
  1616 => x"29b7c449",
  1617 => x"f6e8c191",
  1618 => x"cf4a7481",
  1619 => x"c192c29a",
  1620 => x"70307248",
  1621 => x"72baff4a",
  1622 => x"70986948",
  1623 => x"7487db79",
  1624 => x"29b7c449",
  1625 => x"f6e8c191",
  1626 => x"cf4a7481",
  1627 => x"c392c29a",
  1628 => x"70307248",
  1629 => x"b069484a",
  1630 => x"9d757970",
  1631 => x"87f0c005",
  1632 => x"c848d0ff",
  1633 => x"d4ff78e1",
  1634 => x"c178c548",
  1635 => x"02bfdae7",
  1636 => x"e0c387c3",
  1637 => x"d6e7c178",
  1638 => x"87c602bf",
  1639 => x"c348d4ff",
  1640 => x"d4ff78f0",
  1641 => x"ff0b7b0b",
  1642 => x"e1c848d0",
  1643 => x"78e0c078",
  1644 => x"48dae7c1",
  1645 => x"e7c178c0",
  1646 => x"78c048d6",
  1647 => x"49e2dec2",
  1648 => x"7087f2f9",
  1649 => x"abb7c04b",
  1650 => x"87fefc03",
  1651 => x"4d2648c0",
  1652 => x"4b264c26",
  1653 => x"00004f26",
  1654 => x"00000000",
  1655 => x"711e0000",
  1656 => x"cdfc494a",
  1657 => x"1e4f2687",
  1658 => x"49724ac0",
  1659 => x"e8c191c4",
  1660 => x"79c081f6",
  1661 => x"b7d082c1",
  1662 => x"87ee04aa",
  1663 => x"5e0e4f26",
  1664 => x"0e5d5c5b",
  1665 => x"dcf84d71",
  1666 => x"c44a7587",
  1667 => x"c1922ab7",
  1668 => x"7582f6e8",
  1669 => x"c29ccf4c",
  1670 => x"4b496a94",
  1671 => x"9bc32b74",
  1672 => x"307448c2",
  1673 => x"bcff4c70",
  1674 => x"98714874",
  1675 => x"ecf77a70",
  1676 => x"fe487387",
  1677 => x"000087d8",
  1678 => x"00000000",
  1679 => x"00000000",
  1680 => x"00000000",
  1681 => x"00000000",
  1682 => x"00000000",
  1683 => x"00000000",
  1684 => x"00000000",
  1685 => x"00000000",
  1686 => x"00000000",
  1687 => x"00000000",
  1688 => x"00000000",
  1689 => x"00000000",
  1690 => x"00000000",
  1691 => x"00000000",
  1692 => x"00000000",
  1693 => x"ff1e0000",
  1694 => x"e1c848d0",
  1695 => x"ff487178",
  1696 => x"c47808d4",
  1697 => x"d4ff4866",
  1698 => x"4f267808",
  1699 => x"c44a711e",
  1700 => x"721e4966",
  1701 => x"87deff49",
  1702 => x"c048d0ff",
  1703 => x"262678e0",
  1704 => x"1e731e4f",
  1705 => x"66c84b71",
  1706 => x"4a731e49",
  1707 => x"49a2e0c1",
  1708 => x"2687d9ff",
  1709 => x"4d2687c4",
  1710 => x"4b264c26",
  1711 => x"ff1e4f26",
  1712 => x"ffc34ad4",
  1713 => x"48d0ff7a",
  1714 => x"de78e1c0",
  1715 => x"ecdec27a",
  1716 => x"48497abf",
  1717 => x"7a7028c8",
  1718 => x"28d04871",
  1719 => x"48717a70",
  1720 => x"7a7028d8",
  1721 => x"c048d0ff",
  1722 => x"4f2678e0",
  1723 => x"48d0ff1e",
  1724 => x"7178c9c8",
  1725 => x"08d4ff48",
  1726 => x"1e4f2678",
  1727 => x"eb494a71",
  1728 => x"48d0ff87",
  1729 => x"4f2678c8",
  1730 => x"711e731e",
  1731 => x"fcdec24b",
  1732 => x"87c302bf",
  1733 => x"ff87ebc2",
  1734 => x"c9c848d0",
  1735 => x"c0487378",
  1736 => x"d4ffb0e0",
  1737 => x"dec27808",
  1738 => x"78c048f0",
  1739 => x"c50266c8",
  1740 => x"49ffc387",
  1741 => x"49c087c2",
  1742 => x"59f8dec2",
  1743 => x"c60266cc",
  1744 => x"d5d5c587",
  1745 => x"cf87c44a",
  1746 => x"c24affff",
  1747 => x"c25afcde",
  1748 => x"c148fcde",
  1749 => x"2687c478",
  1750 => x"264c264d",
  1751 => x"0e4f264b",
  1752 => x"5d5c5b5e",
  1753 => x"c24a710e",
  1754 => x"4cbff8de",
  1755 => x"cb029a72",
  1756 => x"91c84987",
  1757 => x"4bfeebc1",
  1758 => x"87c48371",
  1759 => x"4bfeefc1",
  1760 => x"49134dc0",
  1761 => x"dec29974",
  1762 => x"7148bff4",
  1763 => x"08d4ffb8",
  1764 => x"2cb7c178",
  1765 => x"adb7c885",
  1766 => x"c287e704",
  1767 => x"48bff0de",
  1768 => x"dec280c8",
  1769 => x"eefe58f4",
  1770 => x"1e731e87",
  1771 => x"4a134b71",
  1772 => x"87cb029a",
  1773 => x"e6fe4972",
  1774 => x"9a4a1387",
  1775 => x"fe87f505",
  1776 => x"c21e87d9",
  1777 => x"49bff0de",
  1778 => x"48f0dec2",
  1779 => x"c478a1c1",
  1780 => x"03a9b7c0",
  1781 => x"d4ff87db",
  1782 => x"f4dec248",
  1783 => x"dec278bf",
  1784 => x"c249bff0",
  1785 => x"c148f0de",
  1786 => x"c0c478a1",
  1787 => x"e504a9b7",
  1788 => x"48d0ff87",
  1789 => x"dec278c8",
  1790 => x"78c048fc",
  1791 => x"00004f26",
  1792 => x"00000000",
  1793 => x"00000000",
  1794 => x"005f5f00",
  1795 => x"03000000",
  1796 => x"03030003",
  1797 => x"7f140000",
  1798 => x"7f7f147f",
  1799 => x"24000014",
  1800 => x"3a6b6b2e",
  1801 => x"6a4c0012",
  1802 => x"566c1836",
  1803 => x"7e300032",
  1804 => x"3a77594f",
  1805 => x"00004068",
  1806 => x"00030704",
  1807 => x"00000000",
  1808 => x"41633e1c",
  1809 => x"00000000",
  1810 => x"1c3e6341",
  1811 => x"2a080000",
  1812 => x"3e1c1c3e",
  1813 => x"0800082a",
  1814 => x"083e3e08",
  1815 => x"00000008",
  1816 => x"0060e080",
  1817 => x"08000000",
  1818 => x"08080808",
  1819 => x"00000008",
  1820 => x"00606000",
  1821 => x"60400000",
  1822 => x"060c1830",
  1823 => x"3e000103",
  1824 => x"7f4d597f",
  1825 => x"0400003e",
  1826 => x"007f7f06",
  1827 => x"42000000",
  1828 => x"4f597163",
  1829 => x"22000046",
  1830 => x"7f494963",
  1831 => x"1c180036",
  1832 => x"7f7f1316",
  1833 => x"27000010",
  1834 => x"7d454567",
  1835 => x"3c000039",
  1836 => x"79494b7e",
  1837 => x"01000030",
  1838 => x"0f797101",
  1839 => x"36000007",
  1840 => x"7f49497f",
  1841 => x"06000036",
  1842 => x"3f69494f",
  1843 => x"0000001e",
  1844 => x"00666600",
  1845 => x"00000000",
  1846 => x"0066e680",
  1847 => x"08000000",
  1848 => x"22141408",
  1849 => x"14000022",
  1850 => x"14141414",
  1851 => x"22000014",
  1852 => x"08141422",
  1853 => x"02000008",
  1854 => x"0f595103",
  1855 => x"7f3e0006",
  1856 => x"1f555d41",
  1857 => x"7e00001e",
  1858 => x"7f09097f",
  1859 => x"7f00007e",
  1860 => x"7f49497f",
  1861 => x"1c000036",
  1862 => x"4141633e",
  1863 => x"7f000041",
  1864 => x"3e63417f",
  1865 => x"7f00001c",
  1866 => x"4149497f",
  1867 => x"7f000041",
  1868 => x"0109097f",
  1869 => x"3e000001",
  1870 => x"7b49417f",
  1871 => x"7f00007a",
  1872 => x"7f08087f",
  1873 => x"0000007f",
  1874 => x"417f7f41",
  1875 => x"20000000",
  1876 => x"7f404060",
  1877 => x"7f7f003f",
  1878 => x"63361c08",
  1879 => x"7f000041",
  1880 => x"4040407f",
  1881 => x"7f7f0040",
  1882 => x"7f060c06",
  1883 => x"7f7f007f",
  1884 => x"7f180c06",
  1885 => x"3e00007f",
  1886 => x"7f41417f",
  1887 => x"7f00003e",
  1888 => x"0f09097f",
  1889 => x"7f3e0006",
  1890 => x"7e7f6141",
  1891 => x"7f000040",
  1892 => x"7f19097f",
  1893 => x"26000066",
  1894 => x"7b594d6f",
  1895 => x"01000032",
  1896 => x"017f7f01",
  1897 => x"3f000001",
  1898 => x"7f40407f",
  1899 => x"0f00003f",
  1900 => x"3f70703f",
  1901 => x"7f7f000f",
  1902 => x"7f301830",
  1903 => x"6341007f",
  1904 => x"361c1c36",
  1905 => x"03014163",
  1906 => x"067c7c06",
  1907 => x"71610103",
  1908 => x"43474d59",
  1909 => x"00000041",
  1910 => x"41417f7f",
  1911 => x"03010000",
  1912 => x"30180c06",
  1913 => x"00004060",
  1914 => x"7f7f4141",
  1915 => x"0c080000",
  1916 => x"0c060306",
  1917 => x"80800008",
  1918 => x"80808080",
  1919 => x"00000080",
  1920 => x"04070300",
  1921 => x"20000000",
  1922 => x"7c545474",
  1923 => x"7f000078",
  1924 => x"7c44447f",
  1925 => x"38000038",
  1926 => x"4444447c",
  1927 => x"38000000",
  1928 => x"7f44447c",
  1929 => x"3800007f",
  1930 => x"5c54547c",
  1931 => x"04000018",
  1932 => x"05057f7e",
  1933 => x"18000000",
  1934 => x"fca4a4bc",
  1935 => x"7f00007c",
  1936 => x"7c04047f",
  1937 => x"00000078",
  1938 => x"407d3d00",
  1939 => x"80000000",
  1940 => x"7dfd8080",
  1941 => x"7f000000",
  1942 => x"6c38107f",
  1943 => x"00000044",
  1944 => x"407f3f00",
  1945 => x"7c7c0000",
  1946 => x"7c0c180c",
  1947 => x"7c000078",
  1948 => x"7c04047c",
  1949 => x"38000078",
  1950 => x"7c44447c",
  1951 => x"fc000038",
  1952 => x"3c2424fc",
  1953 => x"18000018",
  1954 => x"fc24243c",
  1955 => x"7c0000fc",
  1956 => x"0c04047c",
  1957 => x"48000008",
  1958 => x"7454545c",
  1959 => x"04000020",
  1960 => x"44447f3f",
  1961 => x"3c000000",
  1962 => x"7c40407c",
  1963 => x"1c00007c",
  1964 => x"3c60603c",
  1965 => x"7c3c001c",
  1966 => x"7c603060",
  1967 => x"6c44003c",
  1968 => x"6c381038",
  1969 => x"1c000044",
  1970 => x"3c60e0bc",
  1971 => x"4400001c",
  1972 => x"4c5c7464",
  1973 => x"08000044",
  1974 => x"41773e08",
  1975 => x"00000041",
  1976 => x"007f7f00",
  1977 => x"41000000",
  1978 => x"083e7741",
  1979 => x"01020008",
  1980 => x"02020301",
  1981 => x"7f7f0001",
  1982 => x"7f7f7f7f",
  1983 => x"0808007f",
  1984 => x"3e3e1c1c",
  1985 => x"7f7f7f7f",
  1986 => x"1c1c3e3e",
  1987 => x"10000808",
  1988 => x"187c7c18",
  1989 => x"10000010",
  1990 => x"307c7c30",
  1991 => x"30100010",
  1992 => x"1e786060",
  1993 => x"66420006",
  1994 => x"663c183c",
  1995 => x"38780042",
  1996 => x"6cc6c26a",
  1997 => x"00600038",
  1998 => x"00006000",
  1999 => x"5e0e0060",
  2000 => x"0e5d5c5b",
  2001 => x"c24c711e",
  2002 => x"4dbfcddf",
  2003 => x"1ec04bc0",
  2004 => x"c702ab74",
  2005 => x"48a6c487",
  2006 => x"87c578c0",
  2007 => x"c148a6c4",
  2008 => x"1e66c478",
  2009 => x"dfee4973",
  2010 => x"c086c887",
  2011 => x"eeef49e0",
  2012 => x"4aa5c487",
  2013 => x"f0f0496a",
  2014 => x"87c6f187",
  2015 => x"83c185cb",
  2016 => x"04abb7c8",
  2017 => x"2687c7ff",
  2018 => x"4c264d26",
  2019 => x"4f264b26",
  2020 => x"c24a711e",
  2021 => x"c25ad1df",
  2022 => x"c748d1df",
  2023 => x"ddfe4978",
  2024 => x"1e4f2687",
  2025 => x"4a711e73",
  2026 => x"03aab7c0",
  2027 => x"ccc287d3",
  2028 => x"c405bfdf",
  2029 => x"c24bc187",
  2030 => x"c24bc087",
  2031 => x"c45be3cc",
  2032 => x"e3ccc287",
  2033 => x"dfccc25a",
  2034 => x"9ac14abf",
  2035 => x"49a2c0c1",
  2036 => x"fc87e8ec",
  2037 => x"dfccc248",
  2038 => x"effe78bf",
  2039 => x"4a711e87",
  2040 => x"721e66c4",
  2041 => x"87f9ea49",
  2042 => x"1e4f2626",
  2043 => x"c348d4ff",
  2044 => x"d0ff78ff",
  2045 => x"78e1c048",
  2046 => x"c148d4ff",
  2047 => x"c4487178",
  2048 => x"08d4ff30",
  2049 => x"48d0ff78",
  2050 => x"2678e0c0",
  2051 => x"ccc21e4f",
  2052 => x"e749bfdf",
  2053 => x"dfc287c8",
  2054 => x"bfe848c5",
  2055 => x"c1dfc278",
  2056 => x"78bfec48",
  2057 => x"bfc5dfc2",
  2058 => x"ffc3494a",
  2059 => x"2ab7c899",
  2060 => x"b0714872",
  2061 => x"58cddfc2",
  2062 => x"5e0e4f26",
  2063 => x"0e5d5c5b",
  2064 => x"c8ff4b71",
  2065 => x"c0dfc287",
  2066 => x"7350c048",
  2067 => x"87eee649",
  2068 => x"c24c4970",
  2069 => x"49eecb9c",
  2070 => x"7087cccb",
  2071 => x"c0dfc24d",
  2072 => x"c105bf97",
  2073 => x"66d087e2",
  2074 => x"c9dfc249",
  2075 => x"d60599bf",
  2076 => x"4966d487",
  2077 => x"bfc1dfc2",
  2078 => x"87cb0599",
  2079 => x"fde54973",
  2080 => x"02987087",
  2081 => x"c187c1c1",
  2082 => x"87c1fe4c",
  2083 => x"e2ca4975",
  2084 => x"02987087",
  2085 => x"dfc287c6",
  2086 => x"50c148c0",
  2087 => x"97c0dfc2",
  2088 => x"e3c005bf",
  2089 => x"c9dfc287",
  2090 => x"66d049bf",
  2091 => x"d6ff0599",
  2092 => x"c1dfc287",
  2093 => x"66d449bf",
  2094 => x"caff0599",
  2095 => x"e4497387",
  2096 => x"987087fc",
  2097 => x"87fffe05",
  2098 => x"fbfa4874",
  2099 => x"5b5e0e87",
  2100 => x"f80e5d5c",
  2101 => x"4c4dc086",
  2102 => x"c47ebfec",
  2103 => x"dfc248a6",
  2104 => x"c178bfcd",
  2105 => x"c71ec01e",
  2106 => x"87cefd49",
  2107 => x"987086c8",
  2108 => x"ff87cd02",
  2109 => x"87ebfa49",
  2110 => x"e449dac1",
  2111 => x"4dc187c0",
  2112 => x"97c0dfc2",
  2113 => x"87cf02bf",
  2114 => x"bfd7ccc2",
  2115 => x"c2b9c149",
  2116 => x"7159dbcc",
  2117 => x"c287d4fb",
  2118 => x"4bbfc5df",
  2119 => x"bfdfccc2",
  2120 => x"87e9c005",
  2121 => x"e349fdc3",
  2122 => x"fac387d4",
  2123 => x"87cee349",
  2124 => x"ffc34973",
  2125 => x"c01e7199",
  2126 => x"87e1fa49",
  2127 => x"b7c84973",
  2128 => x"c11e7129",
  2129 => x"87d5fa49",
  2130 => x"f4c586c8",
  2131 => x"c9dfc287",
  2132 => x"029b4bbf",
  2133 => x"ccc287dd",
  2134 => x"c749bfdb",
  2135 => x"987087d5",
  2136 => x"c087c405",
  2137 => x"c287d24b",
  2138 => x"fac649e0",
  2139 => x"dfccc287",
  2140 => x"c287c658",
  2141 => x"c048dbcc",
  2142 => x"c2497378",
  2143 => x"87cd0599",
  2144 => x"e149ebc3",
  2145 => x"497087f8",
  2146 => x"c20299c2",
  2147 => x"734cfb87",
  2148 => x"0599c149",
  2149 => x"f4c387cd",
  2150 => x"87e2e149",
  2151 => x"99c24970",
  2152 => x"fa87c202",
  2153 => x"c849734c",
  2154 => x"87cd0599",
  2155 => x"e149f5c3",
  2156 => x"497087cc",
  2157 => x"d50299c2",
  2158 => x"d1dfc287",
  2159 => x"87ca02bf",
  2160 => x"c288c148",
  2161 => x"c058d5df",
  2162 => x"4cff87c2",
  2163 => x"49734dc1",
  2164 => x"cd0599c4",
  2165 => x"49f2c387",
  2166 => x"7087e3e0",
  2167 => x"0299c249",
  2168 => x"dfc287dc",
  2169 => x"487ebfd1",
  2170 => x"03a8b7c7",
  2171 => x"6e87cbc0",
  2172 => x"c280c148",
  2173 => x"c058d5df",
  2174 => x"4cfe87c2",
  2175 => x"fdc34dc1",
  2176 => x"f9dfff49",
  2177 => x"c2497087",
  2178 => x"87d50299",
  2179 => x"bfd1dfc2",
  2180 => x"87c9c002",
  2181 => x"48d1dfc2",
  2182 => x"c2c078c0",
  2183 => x"c14cfd87",
  2184 => x"49fac34d",
  2185 => x"87d6dfff",
  2186 => x"99c24970",
  2187 => x"87d9c002",
  2188 => x"bfd1dfc2",
  2189 => x"a8b7c748",
  2190 => x"87c9c003",
  2191 => x"48d1dfc2",
  2192 => x"c2c078c7",
  2193 => x"c14cfc87",
  2194 => x"acb7c04d",
  2195 => x"87d3c003",
  2196 => x"c14866c4",
  2197 => x"7e7080d8",
  2198 => x"c002bf6e",
  2199 => x"744b87c5",
  2200 => x"c00f7349",
  2201 => x"1ef0c31e",
  2202 => x"f749dac1",
  2203 => x"86c887cc",
  2204 => x"c0029870",
  2205 => x"dfc287d8",
  2206 => x"6e7ebfd1",
  2207 => x"c491cb49",
  2208 => x"82714a66",
  2209 => x"c5c0026a",
  2210 => x"496e4b87",
  2211 => x"9d750f73",
  2212 => x"87c8c002",
  2213 => x"bfd1dfc2",
  2214 => x"87e2f249",
  2215 => x"bfe3ccc2",
  2216 => x"87ddc002",
  2217 => x"87cbc249",
  2218 => x"c0029870",
  2219 => x"dfc287d3",
  2220 => x"f249bfd1",
  2221 => x"49c087c8",
  2222 => x"c287e8f3",
  2223 => x"c048e3cc",
  2224 => x"f38ef878",
  2225 => x"5e0e87c2",
  2226 => x"0e5d5c5b",
  2227 => x"c24c711e",
  2228 => x"49bfcddf",
  2229 => x"4da1cdc1",
  2230 => x"6981d1c1",
  2231 => x"029c747e",
  2232 => x"a5c487cf",
  2233 => x"c27b744b",
  2234 => x"49bfcddf",
  2235 => x"6e87e1f2",
  2236 => x"059c747b",
  2237 => x"4bc087c4",
  2238 => x"4bc187c2",
  2239 => x"e2f24973",
  2240 => x"0266d487",
  2241 => x"de4987c7",
  2242 => x"c24a7087",
  2243 => x"c24ac087",
  2244 => x"265ae7cc",
  2245 => x"0087f1f1",
  2246 => x"00000000",
  2247 => x"00000000",
  2248 => x"00000000",
  2249 => x"1e000000",
  2250 => x"c8ff4a71",
  2251 => x"a17249bf",
  2252 => x"1e4f2648",
  2253 => x"89bfc8ff",
  2254 => x"c0c0c0fe",
  2255 => x"01a9c0c0",
  2256 => x"4ac087c4",
  2257 => x"4ac187c2",
  2258 => x"4f264872",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
